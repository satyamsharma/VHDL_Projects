Library ieee;
use ieee.std_logic_1164.all;

entity sharma_integration is
port(
in1,in2: in std_logic_vector(7 downto 0);
op: in std_logic_vector(3 downto 0);
start: in std_logic;

result: out std_logic_vector(7 downto 0);
cout, overflow: out std_logic;

--BCD
out1LED,out2LED: out std_logic_vector(7 downto 0);
seg3, seg2, seg1, seg0 : out std_logic_vector(6 downto 0) := "1111111";

signbutton: in std_logic
 );
end sharma_integration;


architecture arch of sharma_integration is
--declare signals in1, in2, out1

  component sharma_eightBitAddSub is
  port(
    a, b : in std_logic_vector(7 downto 0);
    subtract : in std_logic;
    cin : in std_logic;
    cout : out std_logic;
    overflow : out std_logic;
    sum : out std_logic_vector(7 downto 0));
  end component; 

  
  
signal one: std_logic_vector(6 downto 0);
signal ten: std_logic_vector(6 downto 0);
signal hun: std_logic_vector(6 downto 0);
signal sum: std_logic_vector(7 downto 0);
signal sign: std_logic := '0';
signal addsum: std_logic_vector(7 downto 0);
signal couttmp, ovrflotmp : std_logic;

  
  
  
begin
 
process (signbutton)
  begin
    if(signbutton = '0') then
    sign <= not sign;
  end if;
end process;

 
RPPL8 : sharma_eightBitAddSub port map(in1, in2, op(3), op(2), couttmp, ovrflotmp, addsum); 
 
out1LED <= in1;

result <= sum;

process( start )
begin
  if( start = '0') then
    case op is
      when "0011" => --NOTsum
        sum <= not(in1);
		  cout <= '0';
		  overflow <= '0';
      when "0111" => -- OR
        sum <= in1 or in2;
		  cout <= '0';
		  overflow <= '0';
      when "1011" => -- XOR
        sum <= in1 xor in2;
		  cout <= '0';
		  overflow <= '0';
      when "1111" => -- AND
        sum <= in1 and in2;
		  cout <= '0';
		  overflow <= '0';
      when "0001" => -- Left Rotate
        sum <= to_stdlogicvector(to_bitvector(in1) rol 1);
		  cout <= '0';
		  overflow <= '0';
      when "0101" => -- Shift Right
        sum <= to_stdlogicvector(to_bitvector(in1) srl 1);
		  cout <= '0';
		  overflow <= '0';
      when "1001" => -- Shift Left
        sum <= to_stdlogicvector(to_bitvector(in1) sll 1);
		  cout <= '0';
		  overflow <= '0';
      when "1101" => -- Right Rotate
        sum <= to_stdlogicvector(to_bitvector(in1) ror 1);
		  cout <= '0';
		  overflow <= '0';
		when "0010" => -- SLT
			if (to_bitvector(in1) < to_bitvector(in2))
			then sum <= in1;
			elsif (to_bitvector(in1) > to_bitvector(in2))
			then sum <= in2;
			else sum <= "00000000";--(EN = '1') then Q <= D;
			end if;
		when "0110" => -- Add w/ carry
		  sum <= addsum;
		  cout <= couttmp;
		  overflow <= ovrflotmp;
		when "1110" => -- Subtract
		  sum <= addsum;
		  cout <= couttmp;
		  overflow <= ovrflotmp;
		when "1010" => -- Subtract
		  sum <= addsum;
		  cout <= couttmp;
		  overflow <= ovrflotmp;
      when others =>
        NULL;
    end case;
	 	 
	 
  end if;
end process;



seg2 <= hun;
seg1 <= ten;
seg0 <= one;

process(sum, sign) begin
--LOGIC FRIDAY, BCD
if(sign = '0') then
	seg3(0)  <= '1'; 
	one(6) <= ((not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0));
	one(5) <= ((not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0));
	one(4) <= (sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)));
	one(3) <= (sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(1) and sum(0) ) or ( sum(7) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(6)) and sum(5) and sum(4) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(0) ) or ( (not sum(6)) and (not sum(5)) and sum(4) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(4) and sum(3) and sum(2) and sum(0) ) or ( sum(6) and (not sum(5)) and sum(4) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(4) and sum(3) and (not sum(2)) and sum(0) ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(4)) and sum(3) and sum(2) and sum(0) ) or ( sum(6) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(4)) and sum(2) and sum(1) and sum(0));
	one(2) <= (sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(6)) and sum(5) and sum(4) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(0) ) or ( (not sum(6)) and (not sum(5)) and sum(4) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(4) and sum(3) and sum(2) and sum(0) ) or ( sum(6) and (not sum(5)) and sum(4) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(4) and sum(3) and (not sum(2)) and sum(0) ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(5)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(3)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(4)) and sum(3) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(3) and sum(1) and sum(0) ) or ( sum(7) and sum(5) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(5) and (not sum(4)) and (not sum(3)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(3)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(4)) and sum(3) and sum(2) and sum(0) ) or ( (not sum(7)) and (not sum(5)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(3)) and sum(1) and sum(0) ) or ( sum(6) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(4)) and sum(2) and sum(1) and sum(0));
	one(1) <= (sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and (not sum(0)) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and (not sum(0)) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(5)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(3)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(4)) and sum(3) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(3) and sum(1) and sum(0) ) or ( sum(7) and sum(5) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(5) and (not sum(4)) and (not sum(3)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(3)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(5)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(3)) and sum(1) and sum(0));
	one(0) <= (sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and (not sum(1))  ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and sum(2) and (not sum(1))  ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1)  ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and (not sum(1))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and (not sum(1))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and (not sum(2)) and sum(1)  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1))  ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1))  ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1)  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1)  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2)) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and sum(1)  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and sum(1)  ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1))  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2) and (not sum(1))  ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and (not sum(5)) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1))  ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1)  ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1)  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(5)) and sum(4) and sum(3) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(3)) and sum(2) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(1) and sum(0) ) or ( sum(7) and sum(5) and (not sum(4)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and sum(1) and sum(0) ) or ( (not sum(7)) and sum(6) and (not sum(5)) and (not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(3) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(3)) and (not sum(2)) and (not sum(1)) and sum(0) ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(3) and (not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and (not sum(6)) and (not sum(5)) and (not sum(3)) and (not sum(2)) and sum(1) and sum(0));

	ten(6) <= ((not sum(7)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1))  ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(1))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(2)) and sum(1)  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2))  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2)  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2)  ) or ( (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( sum(6) and sum(5) and sum(4) and (not sum(3))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(4)) and sum(3));
	ten(5) <= (sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(2)) and (not sum(1))  ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(1)  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2)  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(1))  ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(2)  ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2))  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and (not sum(3))  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2))  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3))) ;
	ten(4) <= ((not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(1))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(2) and (not sum(1))  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2))  ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(3)) and sum(2)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)));
	ten(3) <= ((not sum(7)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and (not sum(6)) and sum(5) and sum(3) and sum(2) and sum(1)  ) or ( sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1)  ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(1))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(2)) and sum(1)  ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(3)) and (not sum(2))  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(1)  ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(3) and sum(2)  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2)  ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2))  ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2))  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2)  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2)  ) or ( (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and sum(2) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and (not sum(3))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(4)) and sum(3)  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and sum(3));
	ten(2) <= (sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(1)  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2)  ) or ( sum(7) and (not sum(6)) and sum(5) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(2) and sum(1)  ) or ( sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2)) and sum(1)  ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and sum(5) and sum(4) and sum(3) and (not sum(2))  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and (not sum(2)) and (not sum(1))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(1))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(2)) and sum(1)  ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(3)) and (not sum(2))  ) or ( sum(7) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3)  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(1)  ) or ( (not sum(7)) and sum(6) and (not sum(5)) and sum(3) and sum(2)  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(2)) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3)  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2)  ) or ( sum(7) and sum(6) and (not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2))  ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2))  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2)  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2))  ) or ( (not sum(7)) and sum(5) and sum(4) and (not sum(3))  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and sum(2)  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2)  ) or ( (not sum(6)) and (not sum(5)) and sum(4) and (not sum(3)) and (not sum(2))  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and sum(2) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(4)) and (not sum(3))  ) or ( sum(6) and sum(5) and sum(4) and (not sum(3))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(4)) and sum(3)  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and sum(3));
	ten(1) <= (sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(1))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(2) and (not sum(1))  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and (not sum(2)) and (not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and (not sum(3)) and (not sum(2))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and sum(2)  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(2) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(4) and sum(3) and (not sum(2))  ) or ( (not sum(7)) and sum(6) and sum(5) and (not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and sum(3) and sum(2) and sum(1)  ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(3)) and sum(2)  ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(3)) and (not sum(2))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(2)) and sum(1)  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(1)  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(2)) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and (not sum(4)) and sum(3)  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2)  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and sum(3) and (not sum(2))  ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2))  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3)) and sum(2)  ) or ( (not sum(6)) and (not sum(5)) and (not sum(4)) and sum(3) and (not sum(2))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2)  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and sum(2) and sum(1)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(4)) and (not sum(3))  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and sum(3));
	ten(0) <= ((not sum(7)) and sum(6) and sum(5) and (not sum(3)) and sum(2)  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(2))  ) or ( (not sum(7)) and sum(6) and sum(5) and sum(4) and (not sum(3))  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(3)) and (not sum(2))  ) or ( (not sum(7)) and sum(6) and (not sum(4)) and sum(3)  ) or ( sum(6) and (not sum(5)) and (not sum(4)) and sum(3)  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(1)  ) or ( sum(7) and (not sum(6)) and sum(5) and (not sum(4)) and sum(3) and sum(2)  ) or ( sum(7) and (not sum(6)) and sum(5) and sum(4) and (not sum(3)) and (not sum(2))  ) or ( sum(7) and sum(6) and (not sum(5)) and sum(4) and (not sum(3)) and sum(2)  ) or ( (not sum(7)) and (not sum(6)) and (not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and sum(2) and sum(1)  ) or ( (not sum(7)) and (not sum(5)) and (not sum(4)) and sum(3));

	  
	hun(6) <= ((not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( (not sum(6))  ) or ( (not sum(7))) ;
	hun(5) <= ((not sum(7)) and (not sum(4)) and (not sum(3)) and (not sum(2))  ) or ( (not sum(7)) and (not sum(6))  ) or ( (not sum(7)) and (not sum(5))) ;
	hun(4) <= ((not sum(7)) and (not sum(4)) and (not sum(3)) and (not sum(2))  ) or ( sum(7) and sum(6) and sum(5)  ) or ( sum(6) and (not sum(5)) and sum(3)  ) or ( sum(6) and (not sum(5)) and sum(4)  ) or ( (not sum(7)) and (not sum(6))  ) or ( (not sum(7)) and (not sum(5))) ;
	hun(3) <= ((not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( (not sum(6))  ) or ( (not sum(7))) ;
	hun(2) <= ((not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( (not sum(6))  ) or ( (not sum(7))) ;
	hun(1) <= '1';
	hun(0) <= ((not sum(5)) and (not sum(4)) and (not sum(3))  ) or ( (not sum(6))  ) or ( (not sum(7))) ;

else
  
	seg3(0)  <= not sum(7);  
	one(6) <= (sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)));
	one(5) <= (( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1))  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1)  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and sum(1)  ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) );
	one(4) <= (sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)));
	one(3) <= (( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(6) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(6) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(6)) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(0) ) or ( sum(6) and ( not sum(4)) and sum(3) and sum(2) and sum(0) ) or ( ( not sum(6)) and sum(4) and ( not sum(2)) and sum(1) and sum(0) ) or ( sum(6) and ( not sum(4)) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(1)) and sum(0) ) or ( ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and sum(1) and sum(0) ) or ( sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(1)) and sum(0) ) or ( ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and sum(5) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(1) and sum(0));
	one(2) <= (( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(0));
	one(1) <= (sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(1) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and ( not sum(6)) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( sum(7) and ( not sum(6)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and sum(6) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and sum(6) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and sum(4) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and sum(5) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(1)) and sum(0) ) or ( sum(6) and ( not sum(5)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(1) and sum(0) ) or ( ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(1)) and sum(0) ) or ( ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and sum(1) and sum(0) ) or ( sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(1)) and sum(0) ) or ( ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and sum(5) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(1) and sum(0));
	one(0) <= (sum(7) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and sum(1) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and sum(4) and ( not sum(3)) and sum(2) and sum(1) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2)) and ( not sum(1))  ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and sum(2) and ( not sum(1))  ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2) and ( not sum(1))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2)) and sum(1)  ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1)  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1)  ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1)  ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1))  ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1)  ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and sum(5) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(1)) and sum(0) ) or ( sum(6) and ( not sum(5)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(1) and sum(0) ) or ( ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(1)) and sum(0) ) or ( ( not sum(5)) and sum(4) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(3) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and sum(1) and sum(0) ) or ( sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(3)) and sum(2) and ( not sum(1)) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(1)) and sum(0) ) or ( ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(1) and sum(0) ) or ( sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and sum(5) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(1) and sum(0));


	ten(6) <= (sum(7) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3))  ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3))  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(0)) ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(1))  ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and ( not sum(3))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(4)) and sum(3)  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2)) ;
	ten(5) <= (( not sum(6)) and sum(5) and sum(4) and sum(3) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(2)) and ( not sum(1))  ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(2)) and sum(1)  ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(1))  ) or ( ( not sum(6)) and sum(5) and sum(4) and sum(3) and sum(2)  ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2))  ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2)  ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(1))  ) or ( sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and ( not sum(2))  ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3))) ;
	ten(4) <= (sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(2)) and ( not sum(1))  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(2) and ( not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2))  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2)  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2))  ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3)  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and sum(2)  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3))) ;
	ten(3) <= (sum(7) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(3) and sum(2) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2))  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(3) and sum(1)  ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(3) and sum(2)  ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(1)  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3))  ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2)  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3))  ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(2) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(0)) ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(1))  ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and ( not sum(3))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(4)) and sum(3)  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2)  ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(3) );
	ten(2) <= (sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(2) and sum(1) and ( not sum(0)) ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and ( not sum(3)) and sum(2) and sum(0) ) or ( sum(7) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2) and sum(1) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(2)) and sum(1)  ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2))  ) or ( ( not sum(7)) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2)  ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(1))  ) or ( sum(7) and sum(6) and ( not sum(5)) and ( not sum(4)) and sum(3) and ( not sum(2))  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(3)) and ( not sum(2)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(3) and sum(2) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(0) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(1))  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(0)) ) or ( sum(7) and ( not sum(6)) and sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2))  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2)  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(3) and sum(1)  ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(7)) and sum(6) and ( not sum(5)) and sum(3) and sum(2)  ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(1)  ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2)  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and ( not sum(3))  ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(2) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(4)) and ( not sum(3))  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(1))  ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and ( not sum(3))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(4)) and sum(3)  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2)  ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(3)) ;
	ten(1) <= (sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(2) and ( not sum(1)) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(2)) and sum(1) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(2)) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(2) and ( not sum(1))  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and ( not sum(2))  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and ( not sum(3)) and sum(2)  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(4) and sum(3) and ( not sum(2))  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(3)) and ( not sum(2)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(0) ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and sum(3)  ) or ( sum(7) and sum(6) and ( not sum(5)) and sum(4) and sum(3) and sum(2)  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and sum(2)  ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(0)) ) or ( ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3)) and ( not sum(2)) and ( not sum(1))  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(1)  ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2)  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3))  ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(2) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(0)) ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(4)) and ( not sum(3))  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(1))  ) or ( ( not sum(7)) and sum(6) and sum(5) and sum(4) and ( not sum(3))  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2)  ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(3) );
	ten(0) <= (sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(1)) and ( not sum(0)) ) or ( ( not sum(7)) and sum(6) and sum(5) and ( not sum(3)) and sum(2)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(2)) and ( not sum(1)) and sum(0) ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(2))  ) or ( sum(7) and ( not sum(6)) and ( not sum(5)) and sum(4) and ( not sum(3))  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and sum(3) and ( not sum(2)) and ( not sum(0)) ) or ( sum(7) and sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(0) ) or ( ( not sum(7)) and sum(6) and ( not sum(4)) and sum(3)  ) or ( sum(7) and sum(6) and sum(5) and sum(4)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(1)  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and ( not sum(3))  ) or ( sum(6) and sum(5) and ( not sum(4)) and sum(3) and sum(2) and sum(1)  ) or ( sum(7) and ( not sum(6)) and sum(5) and sum(4) and ( not sum(3)) and sum(2)  ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(2) and sum(1)  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(0) ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(1)  ) or ( sum(6) and sum(5) and sum(4) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(7)) and ( not sum(6)) and ( not sum(5)) and ( not sum(3)) and ( not sum(2))  ) or ( ( not sum(6)) and ( not sum(5)) and ( not sum(4)) and sum(3) and sum(2)  ) or ( ( not sum(7)) and ( not sum(5)) and ( not sum(4)) and sum(3) );



	hun(6) <= '1';
	hun(5) <= (( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(0) ) or ( ( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1)  ) or ( sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2))  ) or ( sum(7) and sum(6)  ) or ( ( not sum(6)) and sum(5)  ) or ( ( not sum(7)) and ( not sum(5)) );
	hun(4) <= (( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(0) ) or ( ( not sum(5)) and sum(4) and sum(3) and sum(2) and sum(1)  ) or ( sum(5) and ( not sum(4)) and ( not sum(3)) and ( not sum(2))  ) or ( sum(7) and sum(6)  ) or ( ( not sum(6)) and sum(5)  ) or ( ( not sum(7)) and ( not sum(5)) );
	hun(3) <= '1';
	hun(2) <= '1';
	hun(1) <= '1';
	hun(0) <= '1';
  
  
end if;

end process;

end arch;
